library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ff is
	port(
		clk, rst, mode, pause: in std_logic;
		n0, n1: buffer std_logic_vector(3 downto 0)
	);
end ff;

architecture arc of ff is
	signal cnt: integer := 0;
begin
	process(clk, rst)
	begin
		if (rst = '0') then
			n0 <= "0000";
			n1 <= "0000";
			cnt <= 0;
		elsif (clk'event and clk = '1' and pause = '0') then
			if (mode = '1') then -- clocker (Task#2)
				if (cnt < 4000000) then
					cnt <= cnt + 1;
				else
					cnt <= 0;
				end if;
			end if;
			if (mode = '0' or cnt = 0) then -- +1
				if (n0 = "1001") then
					n0 <= "0000";
					if (n1 = "0101") then
						n1 <= "0000";
					else
						n1 <= n1 + 1;
					end if;
				else
					n0 <= n0 + 1;
				end if;
			end if;
		end if;
	end process;
end arc;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity digit_7 is
	port(
		number: in std_logic_vector(3 downto 0);
		display: out std_logic_vector(6 downto 0)
	);
end digit_7;
architecture arc of digit_7 is
begin
	process(number)
	begin
		case number is
			when "0000"=>display<="1111110";
			when "0001"=>display<="0110000";
			when "0010"=>display<="1101101";
			when "0011"=>display<="1111001";
			when "0100"=>display<="0110011";
			when "0101"=>display<="1011011";
			when "0110"=>display<="0011111";
			when "0111"=>display<="1110000";
			when "1000"=>display<="1111111";
			when "1001"=>display<="1110011";
			when "1010"=>display<="1110111";
			when "1011"=>display<="0011111";
			when "1100"=>display<="1001110";
			when "1101"=>display<="0111101";
			when "1110"=>display<="1001111";
			when "1111"=>display<="1000111";
			when others=>display<="0000000";
		end case;
	end process;
end arc;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity count is
	port(
		clk, rst, mode, pause: in std_logic;
		n0, n1: buffer std_logic_vector(3 downto 0);
		ll, hh: out std_logic_vector(6 downto 0)
	);
end count;

architecture arc of count is
	component ff
		port(
			clk, rst, mode, pause: in std_logic;
			n0, n1: buffer std_logic_vector(3 downto 0)
		);
	end component;
	component digit_7
		port(
			number: in std_logic_vector(3 downto 0);
			display: out std_logic_vector(6 downto 0)
		);	
	end component;
begin
	tmp0: ff port map(clk=>clk, rst=>rst, n0=>n0, n1=>n1, mode=>mode, pause=>pause);
	tmp1: digit_7 port map(number=>n0, display=>ll);
	tmp2: digit_7 port map(number=>n1, display=>hh);
end arc;